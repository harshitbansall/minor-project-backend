* RC Circuit Example
V1 in 0 DC 10
R1 in out 1k
C1 out 0 1uF

.tran 1ms 10ms
.print tran V(out)

.end